module tb;


endmodule