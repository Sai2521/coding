module tt;


endmodule